module APB_SLAVEx(

);

endmodule
